--------------------------------------------------------------------------------
--!
--! @copyright Copyright (c) 2015, DornerWorks Ltd.
--!
--------------------------------------------------------------------------------

library ieee;
use     ieee.std_logic_1164.all;

entity test_axi_gpio is
end entity;

architecture test of test_axi_gpio is
begin
end architecture;
